library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.numeric_std.all;
use std.TEXTIO.ALL ;
 
entity digital_gene is
port (
  reset,clock,start : out std_logic  );
end ;


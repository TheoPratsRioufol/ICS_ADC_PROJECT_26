
wire \vdd3! ;

wire \gnd! ;

wire \vdd! ;

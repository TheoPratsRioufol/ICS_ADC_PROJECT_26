../../digital_part/entity/vhdl.vhd

wire \gnd! ;

wire \vdd! ;
